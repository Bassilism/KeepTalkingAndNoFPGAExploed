----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:56:39 12/14/2020 
-- Design Name: 
-- Module Name:    button_memory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity button_memory is
	port (
			input : in std_logic_vector(3 downto 0)
		);
end button_memory;

architecture Behavioral of button_memory is

begin


end Behavioral;

